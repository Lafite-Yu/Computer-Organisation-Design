`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:11:42 12/13/2017 
// Design Name: 
// Module Name:    MainDec 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MainDec(
	input [31:0] IR_D,
	output [1:0] EXTSrc, 
	output [2:0]Branch, Jump,
	output PCSrc,
	output ALU_BSrc,
	output [3:0] ALUOp,
	output [1:0] MemWrite,
	output [2:0] MemRead,
	output RegWrite,
	output [1:0] RFG_WASrc, GRF_WDSrc, 
	output [2:0] XALU_Op,
	output XALU_Src
    );
	
	`define op IR_D[31:26]
	`define funct IR_D[5:0]
	`define rt IR_D[20:16]
	
	reg [27:0] controls;
	assign {EXTSrc, Branch, Jump, PCSrc, ALU_BSrc, ALUOp, MemWrite, MemRead, RegWrite, RFG_WASrc, GRF_WDSrc, XALU_Op, XALU_Src} = controls;

	always @* begin
		case(`op)
			// Load
			6'b100000: controls = 28'b00_000_000_0_1_0001_00_010_1_00_00_000_0; // lb
			6'b100100: controls = 28'b00_000_000_0_1_0001_00_011_1_00_00_000_0; // lbu
			6'b100001: controls = 28'b00_000_000_0_1_0001_00_100_1_00_00_000_0; // lh
			6'b100101: controls = 28'b00_000_000_0_1_0001_00_101_1_00_00_000_0; // lhu
			6'b100011: controls = 28'b00_000_000_0_1_0001_00_110_1_00_00_000_0; // lw
			// Store
			6'b101000: controls = 28'b00_000_000_0_1_0001_01_000_0_00_00_000_0; // sb
			6'b101001: controls = 28'b00_000_000_0_1_0001_10_000_0_00_00_000_0; // sh
			6'b101011: controls = 28'b00_000_000_0_1_0001_11_000_0_00_00_000_0; // sw
			// R Type
			6'b000000:
				case(`funct)
					// Cal_R
					6'b100000: controls = 28'b00_000_000_0_0_0001_00_000_1_01_01_000_0; // add
					6'b100001: controls = 28'b00_000_000_0_0_0001_00_000_1_01_01_000_0; // addu
					6'b100010: controls = 28'b00_000_000_0_0_0010_00_000_1_01_01_000_0; // sub
					6'b100011: controls = 28'b00_000_000_0_0_0010_00_000_1_01_01_000_0; // subu
					6'b000000: controls = 28'b00_000_000_0_0_0011_00_000_1_01_01_000_0; // sll
					6'b000100: controls = 28'b00_000_000_0_0_0100_00_000_1_01_01_000_0; // sllv
					6'b000010: controls = 28'b00_000_000_0_0_0101_00_000_1_01_01_000_0; // srl
					6'b000110: controls = 28'b00_000_000_0_0_0110_00_000_1_01_01_000_0; // srlv
					6'b000011: controls = 28'b00_000_000_0_0_0111_00_000_1_01_01_000_0; // sra
					6'b000111: controls = 28'b00_000_000_0_0_1000_00_000_1_01_01_000_0; // srav
					6'b100100: controls = 28'b00_000_000_0_0_1001_00_000_1_01_01_000_0; // and
					6'b100101: controls = 28'b00_000_000_0_0_1010_00_000_1_01_01_000_0; // or
					6'b100110: controls = 28'b00_000_000_0_0_1011_00_000_1_01_01_000_0; // xor
					6'b100111: controls = 28'b00_000_000_0_0_1100_00_000_1_01_01_000_0; // nor
					6'b101010: controls = 28'b00_000_000_0_0_1101_00_000_1_01_01_000_0; // slt
					6'b101011: controls = 28'b00_000_000_0_0_1110_00_000_1_01_01_000_0; // sltu
					// Cal_XALU
					6'b010010: controls = 28'b00_000_000_0_0_0000_00_000_1_01_11_001_0; // mflo
					6'b010000: controls = 28'b00_000_000_0_0_0000_00_000_1_01_11_001_1; // mfhi
					6'b010011: controls = 28'b00_000_000_0_0_0000_00_000_0_00_00_010_0; // mtlo
					6'b010001: controls = 28'b00_000_000_0_0_0000_00_000_0_00_00_011_0; // mthi
					6'b011000: controls = 28'b00_000_000_0_0_0000_00_000_0_00_00_110_0; // mult
					6'b011001: controls = 28'b00_000_000_0_0_0000_00_000_0_00_00_111_0; // multu
					6'b011010: controls = 28'b00_000_000_0_0_0000_00_000_0_00_00_100_0; // div
					6'b011011: controls = 28'b00_000_000_0_0_0000_00_000_0_00_00_101_0; // divu
					// Jump
					6'b001001: controls = 28'b00_000_011_1_0_0000_00_000_1_01_10_000_0; // jalr
					6'b001000: controls = 28'b00_000_010_1_0_0000_00_000_0_00_00_000_0; // jr
				endcase
			// Cal_I
			6'b001111: controls = 28'b10_000_000_0_1_0001_00_000_1_00_01_000_0; //lui
			6'b001000: controls = 28'b00_000_000_0_1_0001_00_000_1_00_01_000_0; //addi
			6'b001001: controls = 28'b00_000_000_0_1_0001_00_000_1_00_01_000_0; //addiu
			6'b001100: controls = 28'b01_000_000_0_1_1001_00_000_1_00_01_000_0; //andi
			6'b001101: controls = 28'b01_000_000_0_1_1010_00_000_1_00_01_000_0; //ori
			6'b001110: controls = 28'b01_000_000_0_1_1011_00_000_1_00_01_000_0; //xori
			6'b001010: controls = 28'b00_000_000_0_1_1101_00_000_1_00_01_000_0; //slti
			6'b001011: controls = 28'b00_000_000_0_1_1110_00_000_1_00_01_000_0; //sltiu
			// Branch
			6'b000100: controls = 28'b00_010_000_1_0_0000_00_000_0_00_00_000_0; //beq
			6'b000101: controls = 28'b00_011_000_1_0_0000_00_000_0_00_00_000_0; //bne
			6'b000110: controls = 28'b00_110_000_1_0_0000_00_000_0_00_00_000_0; //blez
			6'b000111: controls = 28'b00_100_000_1_0_0000_00_000_0_00_00_000_0; //bgtz
			6'b000001: 
				case(`rt)
					5'b00000: controls = 28'b00_101_000_1_0_0000_00_000_0_00_00_000_0; //bltz
					5'b00001: controls = 28'b00_111_000_1_0_0000_00_000_0_00_00_000_0; //bgez
				endcase
			// Jump
			6'b000010: controls = 28'b00_000_001_1_0_0000_00_000_0_00_00_000_0; //j
			6'b000011: controls = 28'b00_000_001_1_0_0000_00_000_1_10_10_000_0; //jal
			default: controls = 0;
		endcase
	end
endmodule
